//////////////////////////////////////////////////////////////////////
////                                                              ////
////  can_simple_testbench.v                                      ////
////                                                              ////
////                                                              ////
////  This file is part of the CAN Protocol Controller            ////
////  http://www.opencores.org/projects/can/                      ////
////                                                              ////
////                                                              ////
////  Author(s):                                                  ////
////       Igor Mohor                                             ////
////       igorm@opencores.org                                    ////
////                                                              ////
////                                                              ////
////  All additional information is available in the README.txt   ////
////  file.                                                       ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
////                                                              ////
//// Copyright (C) 2002, 2003 Authors                             ////
////                                                              ////
//// This source file may be used and distributed without         ////
//// restriction provided that this copyright statement is not    ////
//// removed from the file and that any derivative work contains  ////
//// the original copyright notice and the associated disclaimer. ////
////                                                              ////
//// This source file is free software; you can redistribute it   ////
//// and/or modify it under the terms of the GNU Lesser General   ////
//// Public License as published by the Free Software Foundation; ////
//// either version 2.1 of the License, or (at your option) any   ////
//// later version.                                               ////
////                                                              ////
//// This source is distributed in the hope that it will be       ////
//// useful, but WITHOUT ANY WARRANTY; without even the implied   ////
//// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ////
//// PURPOSE.  See the GNU Lesser General Public License for more ////
//// details.                                                     ////
////                                                              ////
//// You should have received a copy of the GNU Lesser General    ////
//// Public License along with this source; if not, download it   ////
//// from http://www.opencores.org/lgpl.shtml                     ////
////                                                              ////
//// The CAN protocol is developed by Robert Bosch GmbH and       ////
//// protected by patents. Anybody who wants to implement this    ////
//// CAN IP core on silicon has to obtain a CAN protocol license  ////
//// from Bosch.                                                  ////
////                                                              ////
//////////////////////////////////////////////////////////////////////


// synopsys translate_off
`include "timescale.v"
// synopsys translate_on
`include "can_defines.v"
`include "can_testbench_defines.v"

module can_simple_testbench();


parameter Tp = 1;
parameter BRP = 2*(`CAN_TIMING0_BRP + 1);


reg         cs_can;
reg         cs_can2;
reg         clk, clk2;
reg         rst;
reg         rx;
wire        tx;
wire        tx_i, tx2_i;
reg         bus_off_on = 1;
reg         bus_off_on2 = 1;
wire        irq;
wire        clkout;

wire        rx_and_tx;

integer     start_tb;
reg   [7:0] tmp_data;
reg         delayed_tx;
reg         tx_bypassed;
reg         extended_mode;

event       igor;

wire [79:0] rx_data, rx_data2;
reg  [63:0] tx_data = 64'h55AA_55AA_55AA_55AA;

reg  tx_start_strobe = 0;
wire tx_succeed, tx_failed;
wire [10:0] id1 = {8'hea, 3'd2};
wire [10:0] id2 = {8'h6a, 3'd2};

can_simple_top i_can_top
(
  .clk_i(clk),
  .rx_i(rx_and_tx),
  .tx_o(tx_i),
  .rst_i(rst),

  .tx_id(id1),
  .tx_data(tx_data),
  .tx_start_strobe(tx_start_strobe),
  .tx_succeed(tx_succeed),
  .tx_failed(tx_failed),
  .rx_data(rx_data),
  .rx_dvalid()
);

// Instantiate can_top module 2
can_simple_top i_can_top2
(
  .clk_i(clk2),
  .rx_i(rx_and_tx),
  .tx_o(tx2_i),
  .rst_i(rst),

  .tx_id(id2),
  .tx_data(tx_data),
  // .tx_start_strobe(tx_start_strobe),
  // .tx_succeed(tx_succeed),
  // .tx_failed(tx_failed),
  .rx_data(rx_data2),
  .rx_dvalid()
);


// Combining tx with the output enable signal.
wire tx_tmp1;
wire tx_tmp2;

assign tx_tmp1 = bus_off_on?  tx_i  : 1'b1;
assign tx_tmp2 = bus_off_on2? tx2_i : 1'b1;

assign tx = tx_tmp1 & tx_tmp2;


// Generate clock signal 25 MHz
// Generate clock signal 16 MHz
initial
begin
  clk=0;
  // forever #20 clk = ~clk;
  // forever #31.25 clk = ~clk; // 16 MHz
  // forever #10.417 clk = ~clk;   // 48 MHz
  forever #8.92857 clk = ~clk;   // 56 MHz
end

initial
begin
  clk2=1;
  forever #28.5 clk2 = ~clk2;
end

initial begin
  rst = 1;
  repeat(5) @(posedge clk);
  rst = 0;
  repeat(50) @(posedge clk);
  @(igor)
 
  @(posedge clk);
  tx_start_strobe = 1;
  @(posedge clk);
  tx_start_strobe = 0;

  wait(tx_succeed | tx_failed);

  repeat(50) @(posedge clk);
  tx_data = 64'h1234_5678_ABCD_EF43;

  @(posedge clk);
  tx_start_strobe = 1;
  @(posedge clk);
  tx_start_strobe = 0;
end

initial
begin
  start_tb = 0;
  cs_can = 0;
  cs_can2 = 0;
  rx = 1;
  extended_mode = 0;
  tx_bypassed = 0;

  repeat(100) @(posedge clk)
  start_tb = 1;
end


// Generating delayed tx signal (CAN transciever delay)
always
begin
  wait (tx);
  repeat (2*BRP) @ (posedge clk);   // 4 time quants delay
  #1 delayed_tx = tx;
  wait (~tx);
  repeat (2*BRP) @ (posedge clk);   // 4 time quants delay
  #1 delayed_tx = tx;
end

//assign rx_and_tx = rx & delayed_tx;   FIX ME !!!
// assign rx_and_tx = /* rx &  */(delayed_tx | tx_bypassed);   // When this signal is on, tx is not looped back to the rx.
assign rx_and_tx = /* rx &  */(tx | tx_bypassed);   // When this signal is on, tx is not looped back to the rx.


// Main testbench
initial
begin
  wait(start_tb);

  #10;
  repeat (1000) @ (posedge clk);
    // Switch-off reset mode

  repeat (BRP) @ (posedge clk);   // At least BRP clocks needed before bus goes to dominant level. Otherwise 1 quant difference is possible
                                  // This difference is resynchronized later.

  // After exiting the reset mode sending bus free
  repeat (11) send_bit(1);

//  test_synchronization;       // test currently switched off
//  test_empty_fifo_ext;        // test currently switched off
//  test_full_fifo_ext;         // test currently switched off
//  send_frame_ext;             // test currently switched off
//  test_empty_fifo;            // test currently switched off
//  test_full_fifo;             // test currently switched off
//  test_reset_mode;              // test currently switched off
//  bus_off_test;               // test currently switched off
//  forced_bus_off;             // test currently switched off
//  send_frame_basic;           // test currently switched on
 send_frame_testBox;
//  send_frame_extended;        // test currently switched off
//  self_reception_request;       // test currently switched off
//  manual_frame_basic;         // test currently switched off
//  manual_frame_ext;           // test currently switched off
//    error_test;
//    register_test;
    // bus_off_recovery_test;

  #1000;
  $display("CAN Testbench finished !");
  $stop;
end


task bus_off_recovery_test;
  begin
    -> igor;

    // Switch-on reset mode



    // Set Clock Divider register
    extended_mode = 1'b1;

    repeat (30) send_bit(1);
    -> igor;
    $display("(%0t) CAN should be idle now", $time);

    // Node 2 sends a message
    // Wait until node 1 receives rx irq

    while (!(tmp_data & 8'h01)) begin

    end

    $display("Frame received by node 1.");

    // Node 1 will send a message and will receive many errors

    fork 
      begin

      end

      begin
        // Waiting until node 1 starts transmitting
        wait (!tx_i);
        repeat (33) send_bit(1);
        repeat (330) send_bit(0);
        repeat (1) send_bit(1);
      end

    join

    // Switch-off reset mode
    repeat (1999) send_bit(1);

    // Switch-on reset mode

    // Switch-off reset mode

    // Wait some time before simulation ends
    repeat (10000) @ (posedge clk);
  end
endtask // bus_off_recovery_test


task error_test;
  begin
    // Switch-off reset mode

    extended_mode = 1'b1;

    repeat (300) send_bit(0);

    $display("Kr neki");

  end
endtask


task register_test;
  integer i, j, tmp;
  begin
    $display("Change mode to extended mode and test registers");
    // Switch-off reset mode



    // Set Clock Divider register
    extended_mode = 1'b1;



    // Switch-off reset mode



    for (i=1; i<128; i=i+1) begin
      for (j=0; j<8; j=j+1) begin


      end
    end

  end
endtask


task send_frame_testBox;    // CAN IP core sends frames
  begin

    ->igor;
  
    fork

      // begin
      //   tx_request_command;
      // end

      // begin
      //   wait (can_simple_testbench.i_can_top.i_can_bsp.go_tx)        // waiting for tx to start
      //   wait (~can_simple_testbench.i_can_top.i_can_bsp.need_to_tx)  // waiting for tx to finish
      //   tx_request_command;                                   // start another tx
      // end

      begin
        // Transmitting acknowledge (for first packet)
        wait (can_simple_testbench.i_can_top.i_can_bsp.tx_state & can_simple_testbench.i_can_top.i_can_bsp.rx_ack & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 0;
        wait (can_simple_testbench.i_can_top.i_can_bsp.rx_ack_lim & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 1;

        // Transmitting acknowledge (for second packet)
        wait (can_simple_testbench.i_can_top.i_can_bsp.tx_state & can_simple_testbench.i_can_top.i_can_bsp.rx_ack & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 0;
        wait (can_simple_testbench.i_can_top.i_can_bsp.rx_ack_lim & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 1;
      end


    join


    #200000;

    // read_receive_buffer2;

    // Read irq register

    #1000;

  end
endtask   // send_frame_testBox


task send_frame_basic;    // CAN IP core sends frames
  begin


    // Enable irqs (basic mode)


    fork

      begin
        #1100;
        $display("\n\nStart receiving data from CAN bus");
        receive_frame(0, 0, {26'h00000e8, 3'h1}, 4'h1, 15'h30bb); // mode, rtr, id, length, crc
        receive_frame(0, 0, {26'h00000e8, 3'h1}, 4'h2, 15'h2da1); // mode, rtr, id, length, crc
        receive_frame(0, 0, {26'h00000ee, 3'h1}, 4'h0, 15'h6cea); // mode, rtr, id, length, crc
        receive_frame(0, 0, {26'h00000e8, 3'h1}, 4'h2, 15'h2da1); // mode, rtr, id, length, crc
        receive_frame(0, 0, {26'h00000ee, 3'h1}, 4'h2, 15'h7b4a); // mode, rtr, id, length, crc
        receive_frame(0, 0, {26'h00000ee, 3'h1}, 4'h1, 15'h00c5); // mode, rtr, id, length, crc
      end

      begin
        // Transmitting acknowledge (for first packet)
        wait (can_simple_testbench.i_can_top.i_can_bsp.tx_state & can_simple_testbench.i_can_top.i_can_bsp.rx_ack & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 0;
        wait (can_simple_testbench.i_can_top.i_can_bsp.rx_ack_lim & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 1;

        // Transmitting acknowledge (for second packet)
        wait (can_simple_testbench.i_can_top.i_can_bsp.tx_state & can_simple_testbench.i_can_top.i_can_bsp.rx_ack & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 0;
        wait (can_simple_testbench.i_can_top.i_can_bsp.rx_ack_lim & can_simple_testbench.i_can_top.i_can_bsp.tx_point);
        #1 rx = 1;
      end


    join

    #200000;

    // read_receive_buffer;

    // Read irq register

    #1000;

  end
endtask   // send_frame_basic

task test_synchronization;
  begin
    // Hard synchronization
    #1 rx=0;
    repeat (2*BRP) @ (posedge clk);
    repeat (8*BRP) @ (posedge clk);
    #1 rx=1;
    repeat (10*BRP) @ (posedge clk);
  
    // Resynchronization on time
    #1 rx=0;
    repeat (10*BRP) @ (posedge clk);
    #1 rx=1;
    repeat (10*BRP) @ (posedge clk);
  
    // Resynchronization late
    repeat (BRP) @ (posedge clk);
    repeat (BRP) @ (posedge clk);
    #1 rx=0;
    repeat (10*BRP) @ (posedge clk);
    #1 rx=1;
  
    // Resynchronization early
    repeat (8*BRP) @ (posedge clk);   // two frames too early
    #1 rx=0;
    repeat (10*BRP) @ (posedge clk);
    #1 rx=1;
    // Resynchronization early
    repeat (11*BRP) @ (posedge clk);   // one frames too late
    #1 rx=0;
    repeat (10*BRP) @ (posedge clk);
    #1 rx=1;

    repeat (10*BRP) @ (posedge clk);
    #1 rx=0;
    repeat (10*BRP) @ (posedge clk);
  end
endtask


task send_bit(logic bit_i);
  integer cnt;
  begin
    #1 rx=bit_i;
    repeat ((`CAN_TIMING1_TSEG1 + `CAN_TIMING1_TSEG2 + 3)*BRP) @ (posedge clk);
  end
endtask


task receive_frame;           // CAN IP core receives frames
  input mode;
  input remote_trans_req;
  input [28:0] id;
  input  [3:0] length;
  input [14:0] crc;

  reg [117:0] data;
  reg         previous_bit;
  reg         stuff;
  reg         tmp;
  reg         arbitration_lost;
  integer     pointer;
  integer     cnt;
  integer     total_bits;
  integer     stuff_cnt;

  begin

    stuff_cnt = 1;
    stuff = 0;

    if(mode)          // Extended format
      data = {id[28:18], 1'b1, 1'b1, id[17:0], remote_trans_req, 2'h0, length};
    else              // Standard format
      data = {id[10:0], remote_trans_req, 1'b0, 1'b0, length};

    if (~remote_trans_req)
      begin
        if(length)    // Send data if length is > 0
          begin
            for (cnt=1; cnt<=(2*length); cnt=cnt+1)  // data   (we are sending nibbles)
              data = {data[113:0], cnt[3:0]};
          end
      end

    // Adding CRC
    data = {data[104:0], crc[14:0]};


    // Calculating pointer that points to the bit that will be send
    if (remote_trans_req)
      begin
        if(mode)          // Extended format
          pointer = 52;
        else              // Standard format
          pointer = 32;
      end
    else
      begin
        if(mode)          // Extended format
          pointer = 52 + 8 * length;
        else              // Standard format
          pointer = 32 + 8 * length;
      end

    // This is how many bits we need to shift
    total_bits = pointer;

    // Waiting until previous msg is finished before sending another one
    if (arbitration_lost)           //  Arbitration lost. Another node is transmitting. We have to wait until it is finished.
      wait ( (~can_simple_testbench.i_can_top.i_can_bsp.error_frame) & 
             (~can_simple_testbench.i_can_top.i_can_bsp.rx_inter   ) & 
             (~can_simple_testbench.i_can_top.i_can_bsp.tx_state   )
           );
    else                            // We were transmitter of the previous frame. No need to wait for another node to finish transmission.
      wait ( (~can_simple_testbench.i_can_top.i_can_bsp.error_frame) & 
             (~can_simple_testbench.i_can_top.i_can_bsp.rx_inter   )
           );
    arbitration_lost = 0;
    
    send_bit(0);                        // SOF
    previous_bit = 0;

    fork 

    begin
      for (cnt=0; cnt<=total_bits; cnt=cnt+1)
        begin
          if (stuff_cnt == 5)
            begin
              stuff_cnt = 1;
              total_bits = total_bits + 1;
              stuff = 1;
              tmp = ~data[pointer+1];
              send_bit(~data[pointer+1]);
              previous_bit = ~data[pointer+1];
            end
          else
            begin
              if (data[pointer] == previous_bit)
                stuff_cnt <= stuff_cnt + 1;
              else
                stuff_cnt <= 1;
              
              stuff = 0;
              tmp = data[pointer];
              send_bit(data[pointer]);
              previous_bit = data[pointer];
              pointer = pointer - 1;
            end
          if (arbitration_lost)
            cnt=total_bits+1;         // Exit the for loop
        end

        // Nothing send after the data (just recessive bit)
        repeat (13) send_bit(1);         // CRC delimiter + ack + ack delimiter + EOF + intermission= 1 + 1 + 1 + 7 + 3
    end

    begin
      while (mode ? (cnt<32) : (cnt<12))
        begin
          #1 wait (can_simple_testbench.i_can_top.sample_point);
          if (mode)
            begin
              if (cnt<32 & tmp & (~rx_and_tx))
                begin
                  arbitration_lost = 1;
                  rx = 1;       // Only recessive is send from now on.
                end
            end
          else
            begin
              if (cnt<12 & tmp & (~rx_and_tx))
                begin
                  arbitration_lost = 1;
                  rx = 1;       // Only recessive is send from now on.
                end
            end
        end
    end

    join

  end
endtask



// State machine monitor (btl)
always @ (posedge clk)
begin
  if(can_simple_testbench.i_can_top.i_can_btl.go_sync & can_simple_testbench.i_can_top.i_can_btl.go_seg1 | can_simple_testbench.i_can_top.i_can_btl.go_sync & can_simple_testbench.i_can_top.i_can_btl.go_seg2 | 
     can_simple_testbench.i_can_top.i_can_btl.go_seg1 & can_simple_testbench.i_can_top.i_can_btl.go_seg2)
    begin
      $display("(%0t) ERROR multiple go_sync, go_seg1 or go_seg2 occurance\n\n", $time);
      #1000;
      $stop;
    end

  if(can_simple_testbench.i_can_top.i_can_btl.sync & can_simple_testbench.i_can_top.i_can_btl.seg1 | can_simple_testbench.i_can_top.i_can_btl.sync & can_simple_testbench.i_can_top.i_can_btl.seg2 | 
     can_simple_testbench.i_can_top.i_can_btl.seg1 & can_simple_testbench.i_can_top.i_can_btl.seg2)
    begin
      $display("(%0t) ERROR multiple sync, seg1 or seg2 occurance\n\n", $time);
      #1000;
      $stop;
    end
end

//
// CRC monitor (used until proper CRC generation is used in testbench
always @ (posedge clk)
begin
  if (can_simple_testbench.i_can_top.i_can_bsp.rx_ack       &
      can_simple_testbench.i_can_top.i_can_bsp.sample_point & 
      can_simple_testbench.i_can_top.i_can_bsp.crc_err
     )
    $display("*E (%0t) ERROR: CRC error (Calculated crc = 0x%0x, crc_in = 0x%0x)", $time, can_simple_testbench.i_can_top.i_can_bsp.calculated_crc, can_simple_testbench.i_can_top.i_can_bsp.crc_in);
end


// form error monitor
always @ (posedge clk)
begin
  if (can_simple_testbench.i_can_top.i_can_bsp.form_err)
    $display("*E (%0t) ERROR: form_error", $time);
end



// acknowledge error monitor
always @ (posedge clk)
begin
  if (can_simple_testbench.i_can_top.i_can_bsp.ack_err)
    $display("*E (%0t) ERROR: acknowledge_error", $time);
end

endmodule

